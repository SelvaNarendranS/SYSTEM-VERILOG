// interface - simple interface using interface in design
// interface
interface intf;
  logic [7:0]a;
  logic [2:0]b;
  logic [7:0]z;
endinterface